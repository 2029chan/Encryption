module kaly_sbox4(x,y);
input [7:0]x;
wire [3:0]i;
wire [3:0]j;
output [7:0] y;
wire [7:0] a[15:0][15:0];

assign j=x[3:0];
assign i=x[7:4];

assign a[0][0]=8'h68;
assign a[0][1]=8'h8d;
assign a[0][2]=8'hca;
assign a[0][3]=8'h4d;
assign a[0][4]=8'h73;
assign a[0][5]=8'h4b;
assign a[0][6]=8'h4e;
assign a[0][7]=8'h2a;
assign a[0][8]=8'hd4;
assign a[0][9]=8'h52;
assign a[0][10]=8'h26;
assign a[0][11]=8'hb3;
assign a[0][12]=8'h54;
assign a[0][13]=8'h1e;
assign a[0][14]=8'h19;
assign a[0][15]=8'h1f;

assign a[1][0]=8'h22;
assign a[1][1]=8'h03;
assign a[1][2]=8'h46;
assign a[1][3]=8'h3d;
assign a[1][4]=8'h2d;
assign a[1][5]=8'h4a;
assign a[1][6]=8'h53;
assign a[1][7]=8'h83;
assign a[1][8]=8'h13;
assign a[1][9]=8'h8a;
assign a[1][10]=8'hb7;
assign a[1][11]=8'hd5;
assign a[1][12]=8'h25;
assign a[1][13]=8'h79;
assign a[1][14]=8'hf5;
assign a[1][15]=8'hbd;

assign a[2][0]=8'h58;
assign a[2][1]=8'h2f;
assign a[2][2]=8'h0d;
assign a[2][3]=8'h02;
assign a[2][4]=8'hed;
assign a[2][5]=8'h51;
assign a[2][6]=8'h9e;
assign a[2][7]=8'h11;
assign a[2][8]=8'hf2;
assign a[2][9]=8'h3e;
assign a[2][10]=8'h55;
assign a[2][11]=8'h5e;
assign a[2][12]=8'hd1;
assign a[2][13]=8'h16;
assign a[2][14]=8'h3c;
assign a[2][15]=8'h66;

assign a[3][0]=8'h70;
assign a[3][1]=8'h5d;
assign a[3][2]=8'hf3;
assign a[3][3]=8'h45;
assign a[3][4]=8'h40;
assign a[3][5]=8'hcc;
assign a[3][6]=8'he8;
assign a[3][7]=8'h94;
assign a[3][8]=8'h56;
assign a[3][9]=8'h08;
assign a[3][10]=8'hce;
assign a[3][11]=8'h1a;
assign a[3][12]=8'h3a;
assign a[3][13]=8'hd2;
assign a[3][14]=8'he1;
assign a[3][15]=8'hdf;

assign a[4][0]=8'hb5;
assign a[4][1]=8'h38;
assign a[4][2]=8'h6e;
assign a[4][3]=8'h0e;
assign a[4][4]=8'he5;
assign a[4][5]=8'hf4;
assign a[4][6]=8'hf9;
assign a[4][7]=8'h86;
assign a[4][8]=8'he9;
assign a[4][9]=8'h4f;
assign a[4][10]=8'hd6;
assign a[4][11]=8'h85;
assign a[4][12]=8'h23;
assign a[4][13]=8'hcf;
assign a[4][14]=8'h32;
assign a[4][15]=8'h99;

assign a[5][0]=8'h31;
assign a[5][1]=8'h14;
assign a[5][2]=8'hae;
assign a[5][3]=8'hee;
assign a[5][4]=8'hc8;
assign a[5][5]=8'h48;
assign a[5][6]=8'hd3;
assign a[5][7]=8'h30;
assign a[5][8]=8'ha1;
assign a[5][9]=8'h92;
assign a[5][10]=8'h41;
assign a[5][11]=8'hb1;
assign a[5][12]=8'h18;
assign a[5][13]=8'hc4;
assign a[5][14]=8'h2c;
assign a[5][15]=8'h71;

assign a[6][0]=8'h72;
assign a[6][1]=8'h44;
assign a[6][2]=8'h15;
assign a[6][3]=8'hfd;
assign a[6][4]=8'h37;
assign a[6][5]=8'hbe;
assign a[6][6]=8'h5f;
assign a[6][7]=8'haa;
assign a[6][8]=8'h9b;
assign a[6][9]=8'h88;
assign a[6][10]=8'hd8;
assign a[6][11]=8'hab;
assign a[6][12]=8'h89;
assign a[6][13]=8'h9c;
assign a[6][14]=8'hfa;
assign a[6][15]=8'h60;

assign a[7][0]=8'hea;
assign a[7][1]=8'hbc;
assign a[7][2]=8'h62;
assign a[7][3]=8'h0c;
assign a[7][4]=8'h24;
assign a[7][5]=8'ha6;
assign a[7][6]=8'ha8;
assign a[7][7]=8'hec;
assign a[7][8]=8'h67;
assign a[7][9]=8'h20;
assign a[7][10]=8'hdb;
assign a[7][11]=8'h7c;
assign a[7][12]=8'h28;
assign a[7][13]=8'hdd;
assign a[7][14]=8'hac;
assign a[7][15]=8'h5b;

assign a[8][0]=8'h34;
assign a[8][1]=8'h7e;
assign a[8][2]=8'h10;
assign a[8][3]=8'hf1;
assign a[8][4]=8'h7b;
assign a[8][5]=8'h8f;
assign a[8][6]=8'h63;
assign a[8][7]=8'ha0;
assign a[8][8]=8'h05;
assign a[8][9]=8'h9a;
assign a[8][10]=8'h43;
assign a[8][11]=8'h77;
assign a[8][12]=8'h21;
assign a[8][13]=8'hbf;
assign a[8][14]=8'h27;
assign a[8][15]=8'h09;

assign a[9][0]=8'hc3;
assign a[9][1]=8'h9f;
assign a[9][2]=8'hb6;
assign a[9][3]=8'hd7;
assign a[9][4]=8'h29;
assign a[9][5]=8'hc2;
assign a[9][6]=8'heb;
assign a[9][7]=8'hc0;
assign a[9][8]=8'ha4;
assign a[9][9]=8'h8b;
assign a[9][10]=8'h8c;
assign a[9][11]=8'h1d;
assign a[9][12]=8'hfb;
assign a[9][13]=8'hff;
assign a[9][14]=8'hc1;
assign a[9][15]=8'hb2;

assign a[10][0]=8'h97;
assign a[10][1]=8'h2e;
assign a[10][2]=8'hf8;
assign a[10][3]=8'h65;
assign a[10][4]=8'hf6;
assign a[10][5]=8'h75;
assign a[10][6]=8'h07;
assign a[10][7]=8'h04;
assign a[10][8]=8'h49;
assign a[10][9]=8'h33;
assign a[10][10]=8'he4;
assign a[10][11]=8'hd9;
assign a[10][12]=8'hb9;
assign a[10][13]=8'hd0;
assign a[10][14]=8'h42;
assign a[10][15]=8'hc7;

assign a[11][0]=8'h6c;
assign a[11][1]=8'h90;
assign a[11][2]=8'h00;
assign a[11][3]=8'h8e;
assign a[11][4]=8'h6f;
assign a[11][5]=8'h50;
assign a[11][6]=8'h01;
assign a[11][7]=8'hc5;
assign a[11][8]=8'hda;
assign a[11][9]=8'h47;
assign a[11][10]=8'h3f;
assign a[11][11]=8'hcd;
assign a[11][12]=8'h69;
assign a[11][13]=8'ha2;
assign a[11][14]=8'he2;
assign a[11][15]=8'h7a;

assign a[12][0]=8'ha7;
assign a[12][1]=8'hc6;
assign a[12][2]=8'h93;
assign a[12][3]=8'h0f;
assign a[12][4]=8'h0a;
assign a[12][5]=8'h06;
assign a[12][6]=8'he6;
assign a[12][7]=8'h2b;
assign a[12][8]=8'h96;
assign a[12][9]=8'ha3;
assign a[12][10]=8'h1c;
assign a[12][11]=8'haf;
assign a[12][12]=8'h6a;
assign a[12][13]=8'h12;
assign a[12][14]=8'h84;
assign a[12][15]=8'h39;

assign a[13][0]=8'he7;
assign a[13][1]=8'hb0;
assign a[13][2]=8'h82;
assign a[13][3]=8'hf7;
assign a[13][4]=8'hfe;
assign a[13][5]=8'h9d;
assign a[13][6]=8'h87;
assign a[13][7]=8'h5c;
assign a[13][8]=8'h81;
assign a[13][9]=8'h35;
assign a[13][10]=8'hde;
assign a[13][11]=8'hb4;
assign a[13][12]=8'ha5;
assign a[13][13]=8'hfc;
assign a[13][14]=8'h80;
assign a[13][15]=8'hef;

assign a[14][0]=8'hcb;
assign a[14][1]=8'hbb;
assign a[14][2]=8'h6b;
assign a[14][3]=8'h76;
assign a[14][4]=8'hba;
assign a[14][5]=8'h5a;
assign a[14][6]=8'h7d;
assign a[14][7]=8'h78;
assign a[14][8]=8'h0b;
assign a[14][9]=8'h95;
assign a[14][10]=8'he3;
assign a[14][11]=8'had;
assign a[14][12]=8'h74;
assign a[14][13]=8'h98;
assign a[14][14]=8'h3b;
assign a[14][15]=8'h36;

assign a[15][0]=8'h64;
assign a[15][1]=8'h6d;
assign a[15][2]=8'hdc;
assign a[15][3]=8'hf0;
assign a[15][4]=8'h59;
assign a[15][5]=8'ha9;
assign a[15][6]=8'h4c;
assign a[15][7]=8'h17;
assign a[15][8]=8'h7f;
assign a[15][9]=8'h91;
assign a[15][10]=8'hb8;
assign a[15][11]=8'hc9;
assign a[15][12]=8'h57;
assign a[15][13]=8'h1b;
assign a[15][14]=8'he0;
assign a[15][15]=8'h61;

assign y=a[i][j];

endmodule

